
module data_modulus(
    input             clk,
    input             rst_n,
    //FFT ST�ӿ�
    input   [23:0]     source_real,   //ʵ�� �з�����
    input   [23:0]     source_imag,   //�鲿 �з�����
    input             source_eop,    //fft����ͨ���������һ�����ݱ�־�ź�
    input             fft_valid,  //�����Ч�źţ�FFT�任��ɺ󣬴��ź��øߣ���ʼ�������
    //ȡģ���������ݽӿ�
    output   [31:0]    fft_data,  //ȡģ�������
    output            data_eop,      //ȡģ���������ֹ�ź�
    output            data_valid     //ȡģ���������Ч�ź�
);

//reg define
reg  [47:0] 	source_data;

wire [47:0]     real_square;
wire [47:0]     image_square;


reg  [23:0]  	data_real;			//ʵ��ԭ��
reg  [23:0]  	data_imag;			//�鲿ԭ��
reg  [7:0]  	source_valid_d;
reg  [7:0] 	    source_eop_d;
wire [31:0]     data_modulus_med;

reg [31:0]    data_modulus;
//*****************************************************
//**                    main code
//***************************************************** 
//wire [9:0] data_modulus_test;
//assign data_modulus_test = fft_data[31:22]; 

assign fft_data = data_modulus ;

assign  data_eop =source_eop;
//assign  data_eop = source_eop_d[7];

  
// �����������ڸ�����Ҫ������Ч�Ķ���ʱ��������  
reg [4:0] counter;  // ʹ��5λ�����������Լ�����17��2^5-1 = 31��  
reg       source_valid;  

always @(posedge clk ) begin  
    if (!rst_n) begin  
        // �첽��λʱ����������������  
        counter <= 5'b0;  
        source_valid <= 1'b0;  
    end else begin  
        // ��⵽a��Чʱ������������  
        if (fft_valid) begin  
            counter <= 5'd17;  // ����Ϊ17���������Ҫ����  
            source_valid <= 1'b1; // �����������Ϊ��Ч  
        end else if (counter > 0) begin  
            // �������ݼ������������Ч  
            counter <= counter - 1'b1;  
            source_valid <= 1'b1;  
        end else begin  
            // ��������0�������Ч  
            source_valid <= 1'b0;  
        end  
    end  
end  
  


/*
//ȡʵ�����鲿��ƽ����
always @ (posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        source_data <= 48'd0;
        data_real   <= 24'd0;
        data_imag   <= 24'd0;
    end
    else begin
        if(source_real[23]==1'b0)               //�ɲ������ԭ��
            data_real <= source_real[23:0];
        else
            data_real <= ~source_real[23:0] + 1'b1;
            
        if(source_imag[23]==1'b0)               //�ɲ������ԭ��
            data_imag <= source_imag[23:0];
        else
            data_imag <= ~source_imag[23:0] + 1'b1;    
                                                //����ԭ��ƽ����
        source_data <= (data_real * data_real) + (data_imag * data_imag);
    end
end
*/

mult_real mult_real (
  .CLK(clk),  // input wire CLK
  .A(source_real),      // input wire A
  .B(source_real),      // input wire B
  .P(real_square)      // output wire P
);

mult_image mult_image (
  .CLK(clk),  // input wire CLK
  .A(source_imag),      // input wire A
  .B(source_imag),      // input wire B
  .P(image_square)      // output wire P
);

//���źŽ��д�����ʱ����
always @ (posedge clk ) begin
    if(!rst_n || !source_valid) begin // 
        source_data <= 48'd0;
    end
    else begin
        source_data <= image_square + real_square;
    end
end

//���źŽ��д�����ʱ����
always @ (posedge clk ) begin
    if(!rst_n) begin
        source_eop_d   <= 8'd0;
        source_valid_d <= 8'd0;
    end
    else begin
        source_valid_d <= {source_valid_d[6:0],source_valid};
        source_eop_d   <= {source_eop_d[6:0],source_eop};
    end
end


always @ (posedge clk ) begin
    if(!rst_n) begin
        data_modulus  <= 32'd0;
    end
    else if(data_valid) begin
        data_modulus<=data_modulus_med[31:9];   //2*data_modulus_med/1024
    end
end


//����cordicģ��,����������
cordic_0 u_cordic_0 (
  .aclk(clk),                                        
  .s_axis_cartesian_tvalid(source_valid),  
  .s_axis_cartesian_tdata(source_data),   
  .m_axis_dout_tvalid(data_valid),         
  .m_axis_dout_tdata(data_modulus_med)            
);

endmodule 
