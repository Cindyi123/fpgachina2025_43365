module fft_test(
    input sys_clk  ,
    input sys_rst_n
    );

wire [31:0]  win_ad_data_out    ;         //�ɼ����adc�������
wire         ad_data_out_en  ;         //�ɼ����adc�������ʹ��

wire [47:0] s_axis_data_tdata;   //fft����ͨ������������
wire        s_axis_data_tvalid;	 //fft����ͨ��������������Чʹ��
wire        s_axis_data_tready;  //fft����ͨ��׼������ź�
wire        s_axis_data_tlast;   //fft����ͨ���������һ�����ݱ�־�ź�
wire        m_axis_data_tvalid;  //fft����ͨ�������������Чʹ��
wire [47:0] m_axis_data_tdata;   //fft����ͨ�����������
wire        m_axis_data_tlast;   //fft����ͨ���������һ�����ݱ�־�ź�
wire [23:0] m_axis_data_tuser;   //fft����ͨ��������ݵ�״̬��Ϣ
wire        fft_eop;             //ȡģ���������ֹ�ź�

    wire          m_axis_data_tvalid_ch3;
     wire  [7 : 0]  m_axis_data_tdata_ch3_med;
     wire  [31 : 0]  m_axis_data_tdata_ch3;
 assign  m_axis_data_tdata_ch3 = m_axis_data_tdata_ch3_med << 16;    


    dds_compiler_0 multi_ch3(
        .aclk(sys_clk),                                // input wire aclk
        .m_axis_data_tvalid(m_axis_data_tvalid_ch3),    // output wire m_axis_data_tvalid
        .m_axis_data_tdata(m_axis_data_tdata_ch3_med),   // output wire [7 : 0] m_axis_data_tdata
        .m_axis_phase_tvalid(),
        .m_axis_phase_tdata()   
    );

//����fifo����ģ�飬adc����
fifo_windows_ctrl u_fifo_ctrl(
	.axi_clk			(sys_clk),         
	.sys_rst_n			(sys_rst_n),              //��λ�źţ��͵�ƽ��Ч

	.ad_clk				(sys_clk),        //��λƫ�ƺ��25mʱ�� 
	.ad_data_in			(m_axis_data_tdata_ch3),            //AD�������� 
    .data_32_en         (m_axis_data_tvalid_ch3),
    
	.s_axis_data_tready	(s_axis_data_tready), //fft����ͨ��׼������ź�
	.s_axis_data_tlast	(s_axis_data_tlast),  //fft����ͨ���������һ�����ݱ�־�ź�

	.win_ad_data_out	(win_ad_data_out),        //�ɼ����adc�������
	.ad_data_out_en     (ad_data_out_en)      //�ɼ����adc�������ʹ��
    
);	
//���ɼ����adc���������Чʹ�ܸ���fft������������Чʹ��
assign  s_axis_data_tvalid =  ad_data_out_en; 
//���ɼ����adc������ݲ�0����fft����������
assign s_axis_data_tdata = {24'b0,win_ad_data_out[23:0]};  

//����fftģ��
xfft_0 xfft_0 (
  .aclk(sys_clk),                             //100mʱ��               
  .aresetn(sys_rst_n),                             //��λ�źţ��͵�ƽ��Ч           
  .s_axis_config_tdata(8'b1),                  //����ͨ�����������ݣ�1��fft   0��ifft
  .s_axis_config_tvalid(1'b1),                 //����ͨ��������������Чʹ��
  .s_axis_config_tready(),                     //�ⲿģ��׼����������ͨ������
  
  .s_axis_data_tdata(s_axis_data_tdata),       //fft����ͨ������������               
  .s_axis_data_tvalid(s_axis_data_tvalid),     //fft����ͨ��������������Чʹ��              
  .s_axis_data_tready(s_axis_data_tready),     //fft����ͨ��׼������ź�          
  .s_axis_data_tlast(s_axis_data_tlast),       //fft����ͨ���������һ�����ݱ�־�ź�           
  
    
  .m_axis_data_tdata(m_axis_data_tdata),       //fft����ͨ�����������              
  .m_axis_data_tuser(m_axis_data_tuser),       //fft����ͨ��������ݵ�״̬��Ϣ              
  .m_axis_data_tvalid(m_axis_data_tvalid),     //fft����ͨ�������������Чʹ��              
  .m_axis_data_tready(1'b1),                   //�ⲿģ��׼����������ͨ������
  .m_axis_data_tlast(m_axis_data_tlast),       //fft����ͨ���������һ�����ݱ�־�ź�               
  
  .m_axis_status_tdata(),                      //fft״̬����ͨ���������
  .m_axis_status_tvalid(),                     //fft״̬����ͨ�����������Чʹ��
  .m_axis_status_tready(1'b1),                 //�ⲿģ��׼������״̬����
  .event_frame_started(),                      
  .event_tlast_unexpected(),         
  .event_tlast_missing(),               
  .event_status_channel_halt(),   
  .event_data_in_channel_halt(), 
  .event_data_out_channel_halt()
);   

 reg [15:0] cnt_fft=16'd0;
 always @(posedge  sys_clk) begin
   if(m_axis_data_tvalid==1)
        cnt_fft<=cnt_fft+1;
    else
        cnt_fft=16'd0;
 end
wire [31:0] fft_data;
wire fft_valid;

//��������ȡģģ��
data_modulus  u_data_modulus(
    .clk					(sys_clk),
    .rst_n					(sys_rst_n),
                     
    .source_real			(m_axis_data_tdata[23:0]),    //ʵ�� �з�����  �������֧������48bits�����ｫ���ݸ�Ϊ1 4 19 ��24λsigned����
    .source_imag			(m_axis_data_tdata[47:24]),  //�鲿 �з�����
    .source_eop				(m_axis_data_tlast),         //fft����ͨ���������һ�����ݱ�־�ź�
    .fft_valid			(m_axis_data_tvalid),        //�����Ч�źţ�FFT�任��ɺ󣬴��ź��øߣ���ʼ�������
    //ȡģ���������ݽӿ�     
    .fft_data		        (fft_data),                  //ȡģ�������
    .data_eop				(fft_eop),                   //ȡģ���������ֹ�ź�
    .data_valid				(fft_valid)                  //ȡģ���������Ч�ź�
);	





endmodule

