

module tb_PID (
    input wire          clk         ,             
    input wire          rst_n       ,           
    input wire [31:0]   P_target    , 
    output reg [31:0]   i_current 
);

// ϵͳ������ʹ�� Q9.23 λ��������ʾ
parameter KE = 32'd4194;    // 0.5e - 3 ת��
parameter TC = 32'd209715200;       // 
parameter A  = 32'd5670699;    // 0.676 ת��Ϊ
parameter B  = 32'd0;         // ϵ�� b
parameter C  = 32'd83886;     // 0.01 ת��Ϊ 
parameter D  = 32'd0;         // ƫ��ϵ�� d

//P_target = 32'd2517;

parameter KP = 32'd41943040;        // ��������
parameter KI = 32'd838861;        // �������棬���ڻ��������С���ɸ���ʵ���������
parameter KD = 32'd83886;        // ΢�����棬����΢�������С���ɸ���ʵ���������

// ʱ�䲽����ʹ�� 23 λ��������ʾ
//parameter TIME_STEP = 23'd8192; // 0.1 ת��Ϊ 23 λ��������
//wire [31:0]   P_target ;
// reg [31:0]   i_current;
// �ڲ�����
wire [31:0] P;
wire [63:0] P_med1,P_med2;             // �⹦��

reg [31:0] error;         // ���
reg [31:0] integral;      // ������
reg [31:0] previous_error; // �ϴ����
reg [31:0] derivative;    // ΢����
reg [31:0] control_signal; // PID ���

// ����⹦��
assign   P_med1 = ((KE * TC) >> 23) + C ;
assign   P_med2 = ((A * i_current) >> 23) + B ;
assign   P = P_med1 * P_med2 >> 23 ;


// PID �������߼�
always @(posedge clk ) begin
    if (!rst_n) begin
        i_current       <= 32'd0;
        error           <= 32'd0;
        integral        <= 32'd0;
        previous_error  <= 32'd0;
        derivative      <= 32'd0;
        control_signal  <= 32'd0;
    end else begin
        // �������
        error <= P_target - P;
        
        // ������
        integral <= integral + error;
        
        // ΢����
        derivative <= error - previous_error ;
        
        // PID ���
        control_signal <= ((KP * error) >> 23) + ((KI * integral) >> 23) + ((KD * derivative) >> 23);
        
        // ������������
        i_current <= i_current + control_signal;
        
        // ���Ƶ�����������
        if (i_current < 32'd0) begin
            i_current <= 32'd0;
        end else if (i_current > 32'd167772 ) begin // ����������Ϊ 20mA
            i_current <= 32'd167772  ;
        end
        
        // �������
        previous_error <= error;
    end
end

endmodule
